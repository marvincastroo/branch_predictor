// Modulo de predictor investigado.

module ();

endmodule